CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
21 1Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 19 80 0 1 11
0 9
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89884e-315 0
0
9 2-In AND~
219 537 44 0 3 22
0 8 5 7
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
391 0 0
2
5.89884e-315 5.26354e-315
0
9 2-In AND~
219 365 35 0 3 22
0 3 4 8
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3124 0 0
2
5.89884e-315 5.30499e-315
0
7 Pulser~
4 44 281 0 10 12
0 18 19 2 20 0 0 5 5 4
8
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3421 0 0
2
5.89884e-315 5.32571e-315
0
2 +V
167 72 52 0 1 3
0 10
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.89884e-315 5.34643e-315
0
6 74112~
219 601 184 0 7 32
0 10 7 2 7 10 21 6
0
0 0 4192 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
5572 0 0
2
5.89884e-315 5.3568e-315
0
6 74112~
219 453 189 0 7 32
0 10 8 2 8 10 22 5
0
0 0 4192 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
8901 0 0
2
5.89884e-315 5.36716e-315
0
6 74112~
219 301 187 0 7 32
0 10 3 2 3 10 23 4
0
0 0 4192 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7361 0 0
2
5.89884e-315 5.37752e-315
0
6 74112~
219 145 187 0 7 32
0 10 9 2 9 10 24 3
0
0 0 4192 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
4747 0 0
2
5.89884e-315 5.38788e-315
0
9 CC 7-Seg~
183 979 230 0 18 19
10 17 16 15 14 13 12 11 2 25
0 0 1 1 1 1 1 1 2
0
0 0 21104 0
7 GREENCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.89884e-315 5.39306e-315
0
6 74LS48
188 852 101 0 14 29
0 6 5 4 3 26 27 11 12 13
14 15 16 17 28
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89884e-315 5.39824e-315
0
37
9 0 0 0 0 0 0 10 0 0 33 4
979 188
982 188
982 151
983 151
0 8 2 0 0 4096 0 0 10 20 0 3
566 272
1000 272
1000 266
4 0 3 0 0 12416 0 11 0 0 16 5
820 92
807 92
807 218
195 218
195 151
3 0 4 0 0 12416 0 11 0 0 13 6
820 83
796 83
796 198
337 198
337 107
325 107
2 0 5 0 0 20608 0 11 0 0 9 6
820 74
784 74
784 175
686 175
686 76
477 76
7 1 6 0 0 4224 0 6 11 0 0 4
625 148
773 148
773 65
820 65
4 0 7 0 0 8192 0 6 0 0 8 3
577 166
558 166
558 146
3 2 7 0 0 4224 0 2 6 0 0 3
558 44
558 148
577 148
7 2 5 0 0 0 0 7 2 0 0 3
477 153
477 53
513 53
4 0 8 0 0 4096 0 7 0 0 11 3
429 171
405 171
405 153
2 0 8 0 0 8192 0 7 0 0 12 3
429 153
404 153
404 35
3 1 8 0 0 4224 0 3 2 0 0 2
386 35
513 35
7 2 4 0 0 0 0 8 3 0 0 3
325 151
325 44
341 44
0 1 3 0 0 0 0 0 3 15 0 3
248 151
248 26
341 26
4 0 3 0 0 0 0 8 0 0 16 3
277 169
248 169
248 151
7 2 3 0 0 0 0 9 8 0 0 2
169 151
277 151
4 0 9 0 0 4224 0 9 0 0 22 3
121 169
18 169
18 148
3 0 2 0 0 0 0 7 0 0 20 2
423 162
423 272
3 0 2 0 0 0 0 8 0 0 20 2
271 160
271 272
3 3 2 0 0 4224 0 4 6 0 0 3
68 272
571 272
571 157
3 3 2 0 0 0 0 4 9 0 0 3
68 272
68 160
115 160
1 2 9 0 0 0 0 1 9 0 0 5
19 92
19 148
18 148
18 151
121 151
5 0 10 0 0 4096 0 7 0 0 30 2
453 201
453 250
5 0 10 0 0 4096 0 8 0 0 30 2
301 199
301 250
5 0 10 0 0 4096 0 6 0 0 30 2
601 196
601 250
1 0 10 0 0 0 0 6 0 0 30 2
601 121
601 91
1 0 10 0 0 0 0 7 0 0 30 2
453 126
453 91
1 0 10 0 0 0 0 8 0 0 30 2
301 124
301 91
1 0 10 0 0 0 0 9 0 0 30 2
145 124
145 91
1 5 10 0 0 8320 0 5 9 0 0 6
72 61
72 91
674 91
674 250
145 250
145 199
7 7 11 0 0 4224 0 11 10 0 0 3
884 65
994 65
994 266
8 6 12 0 0 4224 0 11 10 0 0 3
884 74
988 74
988 266
9 5 13 0 0 4224 0 11 10 0 0 5
884 83
983 83
983 151
982 151
982 266
10 4 14 0 0 4224 0 11 10 0 0 3
884 92
976 92
976 266
11 3 15 0 0 4224 0 11 10 0 0 3
884 101
970 101
970 266
12 2 16 0 0 4224 0 11 10 0 0 3
884 110
964 110
964 266
13 1 17 0 0 4224 0 11 10 0 0 3
884 119
958 119
958 266
2
-16 0 0 0 700 255 0 0 0 3 2 1 18
8 Elephant
0 0 0 21
692 357 913 388
702 365 902 386
21 Christopher Peligrino
-16 0 0 0 700 255 0 0 0 3 2 1 18
8 Elephant
0 0 0 8
694 387 816 418
705 395 804 416
8 BSCpE-1A
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
